3	0.456000	0.388000
3	0.328000	0.480000
3	0.318000	0.646000
3	0.394000	0.774000
3	0.598000	0.844000
4	0.834000	0.708000
3	0.586000	0.494000
3	0.460000	0.474000
3	0.490000	0.652000
3	0.506000	0.802000
4	0.736000	0.772000
3	0.656000	0.574000
4	0.620000	0.656000
3	0.424000	0.572000
4	0.258000	0.586000
4	0.202000	0.786000
3	0.370000	0.890000
3	0.512000	0.902000
3	0.430000	0.696000
3	0.568000	0.772000
4	0.722000	0.908000
3	0.672000	0.778000
3	0.700000	0.692000
4	0.816000	0.832000
4	0.406000	0.280000
4	0.324000	0.336000
4	0.224000	0.514000
4	0.178000	0.656000
3	0.282000	0.770000
3	0.478000	0.550000
3	0.572000	0.602000
4	0.544000	0.318000
4	0.622000	0.396000
4	0.706000	0.488000
4	0.754000	0.564000
4	0.882000	0.738000
4	0.730000	0.926000
4	0.576000	0.940000
4	0.334000	0.954000
4	0.230000	0.884000
4	0.172000	0.528000
4	0.190000	0.442000
4	0.258000	0.382000
4	0.168000	0.608000
4	0.192000	0.732000
