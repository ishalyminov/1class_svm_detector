4	0.460000	0.528000
4	0.430000	0.558000
4	0.444000	0.612000
4	0.530000	0.604000
1	0.490000	0.574000
1	0.520000	0.542000
1	0.506000	0.652000
2	0.132000	0.546000
2	0.214000	0.666000
2	0.330000	0.820000
2	0.598000	0.822000
4	0.582000	0.676000
2	0.588000	0.606000
4	0.514000	0.496000
2	0.340000	0.556000
2	0.308000	0.690000
2	0.372000	0.794000
4	0.430000	0.836000
2	0.598000	0.740000
2	0.506000	0.836000
2	0.414000	0.744000
2	0.510000	0.742000
2	0.560000	0.820000
4	0.472000	0.700000
2	0.386000	0.696000
2	0.346000	0.634000
4	0.390000	0.596000
2	0.308000	0.760000
2	0.392000	0.852000
2	0.246000	0.874000
2	0.046000	0.790000
2	0.150000	0.684000
2	0.262000	0.784000
2	0.294000	0.844000
2	0.254000	0.720000
2	0.262000	0.672000
2	0.170000	0.614000
2	0.048000	0.548000
2	0.072000	0.430000
2	0.146000	0.522000
2	0.226000	0.592000
2	0.290000	0.622000
4	0.332000	0.460000
4	0.382000	0.524000
4	0.436000	0.482000
2	0.592000	0.446000
2	0.664000	0.532000
2	0.564000	0.432000
2	0.438000	0.422000
2	0.262000	0.492000
2	0.726000	0.704000
2	0.858000	0.762000
2	0.670000	0.822000
2	0.762000	0.908000
2	0.500000	0.884000
2	0.632000	0.890000
2	0.644000	0.622000
2	0.810000	0.590000
2	0.686000	0.388000
2	0.514000	0.240000
2	0.616000	0.532000
2	0.694000	0.610000
2	0.800000	0.690000
2	0.472000	0.376000
